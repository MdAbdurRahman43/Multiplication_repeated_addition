`timescale 1ns/1ns
module register_p(y,z,ldp,clrp,clk);
input ldp,clrp,clk;
input [15:0] z;
output [15:0] y;
reg [15:0] out;
assign y=out;
always @(posedge clk)
begin 
if(clrp)
out<=16'h0000;
if(ldp)
out<=z;

end

endmodule
